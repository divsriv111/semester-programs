----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:06:03 05/13/2017 
-- Design Name: 
-- Module Name:    SIPO_shift - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SIPO_shift is
    Port ( clk,si : in  STD_LOGIC;
           po : inout  STD_LOGIC_VECTOR(3 downto 0));
end SIPO_shift;
architecture Behavioral of SIPO_shift is
begin
process(clk)
begin
if(clk'event and clk='1')then
po(3 downto 1)<=po(2 downto 0);
po(0)<=si;
end if;
end process;
end Behavioral;

