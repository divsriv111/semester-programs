----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:37:08 03/15/2018 
-- Design Name: 
-- Module Name:    ex4_q2_1x8DMUX - Structural 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ex4_q2_1x8DMUX is
    Port ( d,e,s0,s1 : in  STD_LOGIC;
           i1,i2,i3,i4,i5,i6,i7,i8 : out  STD_LOGIC);
end ex4_q2_1x8DMUX;

architecture Structural of ex4_q2_1x8DMUX is
component ex4_q2_1x4DMUX
port( d,e,s0,s1 : in std_logic;
		i1,i2,i3,i4 : out std_logic);
end component;
begin
dm1:ex4_q2_1x4DMUX port map(d,NOT e,s0,s1,i1,i2,i3,i4);
dm2:ex4_q2_1x4DMUX port map(d,e,s0,s1,i5,i6,i7,i8);
end Structural;

