----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:12:08 03/14/2018 
-- Design Name: 
-- Module Name:    ex2_q2_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ex2_q2_1 is
    Port ( x,y,a,b : in  STD_LOGIC;
           o : out  STD_LOGIC);
end ex2_q2_1;

architecture Behavioral of ex2_q2_1 is

begin
process(x,y,a,b)
begin

if(x='0' and y='0') then
o <= a AND b;
elsif(x='0' and y='1') then
o <= a OR b;
elsif(x='1' and y='0') then
o <= a NOR b;
else
o <= a NAND b;
end if;

end process;
end Behavioral;

